library IEEE;
use IEEE.std_logic_1164.all;

entity top is
  port (
    clk: in std_logic;
  );
end entity top;
